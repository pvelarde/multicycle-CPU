`timescale 1ns / 1ps

module top_module(clock, reset, alu_output);
input clock;
input reset;
output [31:0] alu_output;




endmodule
